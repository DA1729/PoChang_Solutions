module s_prior_1 (
    input wire [0:11] A,
    output reg [0:3] y
);

always @ *

begin

casez (A)
    12'b1???????????: y = 4'b0000;
    12'b01??????????: y = 4'b0001;
    12'b001?????????: y = 4'b0010;
    12'b0001????????: y = 4'b0011;
    12'b00001???????: y = 4'b0100;
    12'b000001??????: y = 4'b0101;
    12'b0000001?????: y = 4'b0110;
    12'b00000001????: y = 4'b0111;
    12'b000000001???: y = 4'b1000;
    12'b0000000001??: y = 4'b1001;
    12'b00000000001?: y = 4'b1010;
    12'b000000000001: y = 4'b1011;
    default: y = 4'b0000;
endcase
end 

endmodule